/*  # Template matching - Testbench
 *
 *  The template matching testbench will test linebuffer, SAD, and linecounter
 *  module as integrated template matching procedure. The template matching
 *  testbench will load black-and-white source image and the template image
 *  to their apropriate registers.
 */

module bench_template_matching;
